module mux_4x1_trans_tb();
reg a;
reg b;
reg c;
reg d;
reg s1;
reg s2;
wire res;

mux_4x1_trans mux_4x1_trans_tb(
	.d0(a),
	.d1(b),
	.d2(c),
	.d3(d),
	.s0(s1),
	.s1(s2),
	.result(res)
);

	initial
		begin
				s2 = 0; s1 = 0; d = 0; c = 0; b = 0; a = 0; 
			#10 s2 = 0; s1 = 0; d = 0; c = 0; b = 0; a = 1; 
			#10 s2 = 0; s1 = 0; d = 0; c = 0; b = 1; a = 0; 
			#10 s2 = 0; s1 = 0; d = 0; c = 0; b = 1; a = 1; 
			#10 s2 = 0; s1 = 0; d = 0; c = 1; b = 0; a = 0; 
			#10 s2 = 0; s1 = 0; d = 0; c = 1; b = 0; a = 1; 
			#10 s2 = 0; s1 = 0; d = 0; c = 1; b = 1; a = 0; 
			#10 s2 = 0; s1 = 0; d = 0; c = 1; b = 1; a = 1; 
			#10 s2 = 0; s1 = 0; d = 1; c = 0; b = 0; a = 0; 
			#10 s2 = 0; s1 = 0; d = 1; c = 0; b = 0; a = 1; 
			#10 s2 = 0; s1 = 0; d = 1; c = 0; b = 1; a = 0; 
			#10 s2 = 0; s1 = 0; d = 1; c = 0; b = 1; a = 1; 
			#10 s2 = 0; s1 = 0; d = 1; c = 1; b = 0; a = 0; 
			#10 s2 = 0; s1 = 0; d = 1; c = 1; b = 0; a = 1; 
			#10 s2 = 0; s1 = 0; d = 1; c = 1; b = 1; a = 0; 
			#10 s2 = 0; s1 = 0; d = 1; c = 1; b = 1; a = 1; 
			#10 s2 = 0; s1 = 1; d = 0; c = 0; b = 0; a = 0; 
			#10 s2 = 0; s1 = 1; d = 0; c = 0; b = 0; a = 1; 
			#10 s2 = 0; s1 = 1; d = 0; c = 0; b = 1; a = 0; 
			#10 s2 = 0; s1 = 1; d = 0; c = 0; b = 1; a = 1; 
			#10 s2 = 0; s1 = 1; d = 0; c = 1; b = 0; a = 0; 
			#10 s2 = 0; s1 = 1; d = 0; c = 1; b = 0; a = 1; 
			#10 s2 = 0; s1 = 1; d = 0; c = 1; b = 1; a = 0; 
			#10 s2 = 0; s1 = 1; d = 0; c = 1; b = 1; a = 1; 
			#10 s2 = 0; s1 = 1; d = 1; c = 0; b = 0; a = 0; 
			#10 s2 = 0; s1 = 1; d = 1; c = 0; b = 0; a = 1; 
			#10 s2 = 0; s1 = 1; d = 1; c = 0; b = 1; a = 0; 
			#10 s2 = 0; s1 = 1; d = 1; c = 0; b = 1; a = 1; 
			#10 s2 = 0; s1 = 1; d = 1; c = 1; b = 0; a = 0; 
			#10 s2 = 0; s1 = 1; d = 1; c = 1; b = 0; a = 1; 
			#10 s2 = 0; s1 = 1; d = 1; c = 1; b = 1; a = 0; 
			#10 s2 = 0; s1 = 1; d = 1; c = 1; b = 1; a = 1; 
			#10 s2 = 1; s1 = 0; d = 0; c = 0; b = 0; a = 0; 
			#10 s2 = 1; s1 = 0; d = 0; c = 0; b = 0; a = 1; 
			#10 s2 = 1; s1 = 0; d = 0; c = 0; b = 1; a = 0; 
			#10 s2 = 1; s1 = 0; d = 0; c = 0; b = 1; a = 1; 
			#10 s2 = 1; s1 = 0; d = 0; c = 1; b = 0; a = 0; 
			#10 s2 = 1; s1 = 0; d = 0; c = 1; b = 0; a = 1; 
			#10 s2 = 1; s1 = 0; d = 0; c = 1; b = 1; a = 0; 
			#10 s2 = 1; s1 = 0; d = 0; c = 1; b = 1; a = 1; 
			#10 s2 = 1; s1 = 0; d = 1; c = 0; b = 0; a = 0; 
			#10 s2 = 1; s1 = 0; d = 1; c = 0; b = 0; a = 1; 
			#10 s2 = 1; s1 = 0; d = 1; c = 0; b = 1; a = 0; 
			#10 s2 = 1; s1 = 0; d = 1; c = 0; b = 1; a = 1; 
			#10 s2 = 1; s1 = 0; d = 1; c = 1; b = 0; a = 0; 
			#10 s2 = 1; s1 = 0; d = 1; c = 1; b = 0; a = 1; 
			#10 s2 = 1; s1 = 0; d = 1; c = 1; b = 1; a = 0; 
			#10 s2 = 1; s1 = 0; d = 1; c = 1; b = 1; a = 1; 
			#10 s2 = 1; s1 = 1; d = 0; c = 0; b = 0; a = 0; 
			#10 s2 = 1; s1 = 1; d = 0; c = 0; b = 0; a = 1; 
			#10 s2 = 1; s1 = 1; d = 0; c = 0; b = 1; a = 0; 
			#10 s2 = 1; s1 = 1; d = 0; c = 0; b = 1; a = 1; 
			#10 s2 = 1; s1 = 1; d = 0; c = 1; b = 0; a = 0; 
			#10 s2 = 1; s1 = 1; d = 0; c = 1; b = 0; a = 1; 
			#10 s2 = 1; s1 = 1; d = 0; c = 1; b = 1; a = 0; 
			#10 s2 = 1; s1 = 1; d = 0; c = 1; b = 1; a = 1; 
			#10 s2 = 1; s1 = 1; d = 1; c = 0; b = 0; a = 0; 
			#10 s2 = 1; s1 = 1; d = 1; c = 0; b = 0; a = 1; 
			#10 s2 = 1; s1 = 1; d = 1; c = 0; b = 1; a = 0; 
			#10 s2 = 1; s1 = 1; d = 1; c = 0; b = 1; a = 1; 
			#10 s2 = 1; s1 = 1; d = 1; c = 1; b = 0; a = 0; 
			#10 s2 = 1; s1 = 1; d = 1; c = 1; b = 0; a = 1; 
			#10 s2 = 1; s1 = 1; d = 1; c = 1; b = 1; a = 0; 
			#10 s2 = 1; s1 = 1; d = 1; c = 1; b = 1; a = 1; 
		end

	initial
		begin
			$dumpfile("mux_4x1_trans.vcd");
			$dumpvars(0, mux_4x1_trans_tb);
			$monitor("time = %2d, abit = %1b, bbit = %1b, cbit = %1b, dbit = %1b, s1bit = %1b, s2bit = %1b, result = %1b", $time, a, b, c, d, s1, s2, res);
		end

endmodule