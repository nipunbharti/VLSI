module multiplier15bit(input [15:0] a, input [15:0] b, output [31:0] result);

	assign result = a * b;

endmodule