module subtracter32bit(input [31:0] a, input [31:0] b, output [32:0] result);

	assign result = a - b;

endmodule